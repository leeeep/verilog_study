module alu(
);

hehehe;
dssds;
endmodule