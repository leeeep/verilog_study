module alu(
);

hehehe;

endmodule