module alu(
);
